// this is test file for git
module test()
